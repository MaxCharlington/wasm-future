`include "stack.svh"

// Operations
`define INDEX_RESET           4
`define INDEX_RESET_AND_PUSH  5
`define UNDERFLOW_GET         6
`define UNDERFLOW_SET         7

// Errors
`define BAD_OFFSET 3
